LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SEQ_ENCODER IS
	PORT(MSG: IN STD_LOGIC;
		  CLK: IN STD_LOGIC;
		  NRST: IN STD_LOGIC;
		  ENC_MSG: OUT STD_LOGIC);
END SEQ_ENCODER;

ARCHITECTURE STRUCTURAL OF SEQ_ENCODER IS

--SAIDA DOS XORS
SIGNAL S_XOR0 : STD_LOGIC;
SIGNAL S_XOR1 : STD_LOGIC;
SIGNAL S_XOR2 : STD_LOGIC;
SIGNAL S_XOR3 : STD_LOGIC;
--SAIDA DOS REGISTOS
SIGNAL S_REG0 : STD_LOGIC;
SIGNAL S_REG1 : STD_LOGIC;
SIGNAL S_REG2 : STD_LOGIC;
SIGNAL S_REG3 : STD_LOGIC;

--SAIDA DOS ANDS
SIGNAL S_AND0 : STD_LOGIC;
SIGNAL S_AND1 : STD_LOGIC;
SIGNAL S_AND2 : STD_LOGIC;
SIGNAL S_AND3 : STD_LOGIC;

--SAIDA DO 4MUX1
SIGNAL S_MUX4 : STD_LOGIC;

--SAIDA DO 2MUX1
SIGNAL S_MUX2 : STD_LOGIC;

--SINAL CONTROLO DOS ANDS
SIGNAL S_ENP0 : STD_LOGIC;
SIGNAL S_ENP1 : STD_LOGIC;
SIGNAL S_ENP2 : STD_LOGIC;
SIGNAL S_ENP3 : STD_LOGIC;

--SINAL CONTROLO DO 4MUX1
SIGNAL S_CMUX4 : STD_LOGIC_VECTOR(1 DOWNTO 0);

--SINAL CONTROLO DO 2MUX1
SIGNAL S_CMUX2 : STD_LOGIC;

--SAIDA DO CNT4BIT
SIGNAL S_ADDR : STD_LOGIC_VECTOR(3 DOWNTO 0);

--SAIDA DA RAM
SIGNAL S_CTRLB : STD_LOGIC_VECTOR(6 DOWNTO 0); 

BEGIN

	REG0: WORK.FLIPFLOPDSIMUL PORT MAP (CLK,S_XOR0,'1',NRST,S_REG0,OPEN);
	REG1: WORK.FLIPFLOPDSIMUL PORT MAP (CLK,S_XOR1,'1',NRST,S_REG1,OPEN);
	REG2: WORK.FLIPFLOPDSIMUL PORT MAP (CLK,S_XOR2,'1',NRST,S_REG2,OPEN);
	REG3: WORK.FLIPFLOPDSIMUL PORT MAP (CLK,S_XOR3,'1',NRST,S_REG3,OPEN);

	AND0: WORK.AANDB PORT MAP (MSG,S_ENP0,S_AND0);
	AND1: WORK.AANDB PORT MAP (MSG,S_ENP1,S_AND1);
	AND2: WORK.AANDB PORT MAP (MSG,S_ENP2,S_AND2);
	AND3: WORK.AANDB PORT MAP (MSG,S_ENP3,S_AND3);
	
	XOR0: WORK.AXORB PORT MAP (S_AND0,S_REG0,S_XOR0);
	XOR1: WORK.AXORB PORT MAP (S_AND1,S_REG1,S_XOR1);
	XOR2: WORK.AXORB PORT MAP (S_AND2,S_REG2,S_XOR2);
	XOR3: WORK.AXORB PORT MAP (S_AND3,S_REG3,S_XOR3);
	
	MUX4TO1: WORK.MULT4TO1 PORT MAP (S_XOR0,S_XOR1,S_XOR2,S_XOR3,S_CMUX4,S_MUX4);
	
	MUX2TO1: WORK.MULT2TO1 PORT MAP (MSG,S_MUX4,S_CMUX2,ENC_MSG);
	
	CNT0: WORK.COUNTER4BIT PORT MAP (CLK,NRST,S_ADDR,OPEN);
	
	ROM0: WORK.SEQ_ENCODER_CTRL_ROM PORT MAP (S_ADDR,S_CTRLB);
	
	S_ENP0<=S_CTRLB(6);
	S_ENP1<=S_CTRLB(5);
	S_ENP2<=S_CTRLB(4);
	S_ENP3<=S_CTRLB(3);
	S_CMUX2<=S_CTRLB(2);
	S_CMUX4<=S_CTRLB(1)&S_CTRLB(0);
	

END STRUCTURAL;

------------------------
--ROM DE CONTROLO

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY SEQ_ENCODER_CTRL_ROM IS
	PORT(ADDR: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		  CTRLBITS: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END SEQ_ENCODER_CTRL_ROM;

ARCHITECTURE BEHAVIORAL OF SEQ_ENCODER_CTRL_ROM IS

	--S_ENP0,S_ENP1,S_ENP2,S_ENP3,S_CMUX2,S_CMUX4_0,S_CMUX4_1
	TYPE TROM IS ARRAY (0 TO 14) OF STD_LOGIC_VECTOR(6 DOWNTO 0); 
	CONSTANT ROM_TABLE : TROM := (
		"1100000",
		"1010000",
		"1001000",
		"0110000",
		"0101000",
		"0011000",
		"1110000",
		"1101000",
		"1011000",
		"0111000",
		"1111000",
		--PARITY
		"0000100",
		"0000101",
		"0000110",
		"0000111"
		);
BEGIN
		CTRLBITS<=ROM_TABLE(TO_INTEGER(UNSIGNED(ADDR)));
END BEHAVIORAL;
