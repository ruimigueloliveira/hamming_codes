LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PARALLEL_DECODER IS
  PORT( CODED_MESSAGE : IN  STD_LOGIC_VECTOR(14 DOWNTO 0);
		  MESSAGE : OUT STD_LOGIC_VECTOR(10 DOWNTO 0));
END PARALLEL_DECODER;

ARCHITECTURE STRUCTURAL OF PARALLEL_DECODER IS

SIGNAL S_PARITY_BITS : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL S_MASK : STD_LOGIC_VECTOR(10 DOWNTO 0);

BEGIN

	PARITY_BITS: WORK.PARITY_BITS_CALCULATOR PORT MAP(CODED_MESSAGE, S_PARITY_BITS);
	MASK: WORK.DECODER_4TO11 PORT MAP(S_PARITY_BITS, S_MASK);
	
	-- BIT CORRECTION
	MESSAGE(0) <= CODED_MESSAGE(0) XOR S_MASK(0);
	MESSAGE(1) <= CODED_MESSAGE(1) XOR S_MASK(1);
	MESSAGE(2) <= CODED_MESSAGE(2) XOR S_MASK(2);
	MESSAGE(3) <= CODED_MESSAGE(3) XOR S_MASK(3);
	MESSAGE(4) <= CODED_MESSAGE(4) XOR S_MASK(4);
	MESSAGE(5) <= CODED_MESSAGE(5) XOR S_MASK(5);
	MESSAGE(6) <= CODED_MESSAGE(6) XOR S_MASK(6);
	MESSAGE(7) <= CODED_MESSAGE(7) XOR S_MASK(7);
	MESSAGE(8) <= CODED_MESSAGE(8) XOR S_MASK(8);
	MESSAGE(9) <= CODED_MESSAGE(9) XOR S_MASK(9);
	MESSAGE(10) <= CODED_MESSAGE(10) XOR S_MASK(10);
	
END STRUCTURAL;