LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY INC4BIT IS
  PORT (A : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        S : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		  OVERFLOW : OUT STD_LOGIC);
END INC4BIT;

ARCHITECTURE STRUCTURAL OF INC4BIT IS

SIGNAL S_COUT0 : STD_LOGIC;
SIGNAL S_COUT1 : STD_LOGIC;
SIGNAL S_COUT2 : STD_LOGIC;

BEGIN
	HA0: WORK.HALFADDER1BIT PORT MAP (A(0), '1', S(0), S_COUT0);
	HA1: WORK.HALFADDER1BIT PORT MAP (A(1), S_COUT0, S(1), S_COUT1);
	HA2: WORK.HALFADDER1BIT PORT MAP (A(2), S_COUT1, S(2), S_COUT2);
	HA3: WORK.HALFADDER1BIT PORT MAP (A(3), S_COUT2, S(3), OVERFLOW);
END STRUCTURAL;