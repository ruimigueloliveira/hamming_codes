LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MULT2TO1 IS
  PORT (X0, X1: IN STD_LOGIC;
        S: IN STD_LOGIC;
        Y: OUT STD_LOGIC);
END MULT2TO1;

ARCHITECTURE BEHAVIORAL OF MULT2TO1 IS
BEGIN
  Y <= (X0 AND NOT S) OR (X1 AND S);
END BEHAVIORAL;