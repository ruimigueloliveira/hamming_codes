LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY HALFADDER1BIT IS
  PORT (A,B : IN STD_LOGIC;
        S,COUT: OUT STD_LOGIC);
END HALFADDER1BIT;

ARCHITECTURE BEHAVIORAL OF HALFADDER1BIT IS
BEGIN
	S <= A XOR B;
	COUT <= A AND B;
END BEHAVIORAL;