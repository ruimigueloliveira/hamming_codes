LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PARALLEL_ENCODER IS
    PORT ( M01, M02, M03, M04, M05, M06, M07, M08, M09, M10, M11: IN STD_LOGIC;
			  X01, X02, X03, X04, X05, X06, X07, X08, X09, X10, X11, X12, X13, X14, X15: OUT STD_LOGIC );
END PARALLEL_ENCODER;

ARCHITECTURE BEHAVIORAL OF PARALLEL_ENCODER IS

-- LEVEL ONE
SIGNAL XOR_M01_M07, XOR_M08_M11, XOR_M02_M03, XOR_M04_M05, XOR_M06_M09, XOR_M10_M11, XOR_M02_M04, XOR_M03_M05: STD_LOGIC;

-- LEVEL TWO
SIGNAL XOR_M01_M07_M08_M11, XOR_M02_M03_M09, XOR_M04_M05_M10, XOR_M06_M09_M10_M11, XOR_M02_M04_M07, XOR_M03_M05_M08: STD_LOGIC;


BEGIN

	X01 <= M01;
	X02 <= M02;
	X03 <= M03;
	X04 <= M04;
	X05 <= M05;
	X06 <= M06;
	X07 <= M07;
	X08 <= M08;
	X09 <= M09;
	X10 <= M10;
	X11 <= M11;
	
	-- LEVEL ONE
	XOR_M01_M07 <= M01 XOR M07;
	XOR_M08_M11 <= M08 XOR M11;
	XOR_M02_M03 <= M02 XOR M03;
	XOR_M04_M05 <= M04 XOR M05;
	XOR_M06_M09 <= M06 XOR M09;
	XOR_M10_M11 <= M10 XOR M11;
	XOR_M02_M04 <= M02 XOR M04;
	XOR_M03_M05 <= M03 XOR M05;
	
	-- LEVEL TWO
	XOR_M01_M07_M08_M11 <= XOR_M01_M07 XOR XOR_M08_M11;
	XOR_M02_M03_M09 <= XOR_M02_M03 XOR M09;
	XOR_M04_M05_M10 <= XOR_M04_M05 XOR M10;
	XOR_M06_M09_M10_M11 <= XOR_M06_M09 XOR XOR_M10_M11;
	XOR_M02_M04_M07 <= XOR_M02_M04 XOR M07;
	XOR_M03_M05_M08 <= XOR_M03_M05 XOR M08;
	
	-- LEVEL THREE
	X12 <= XOR_M01_M07_M08_M11 XOR XOR_M02_M03_M09; 
	X13 <= XOR_M01_M07_M08_M11 XOR XOR_M04_M05_M10; 
	X14 <= XOR_M06_M09_M10_M11 XOR XOR_M02_M04_M07; 
	X15 <= XOR_M06_M09_M10_M11 XOR XOR_M03_M05_M08; 
	
END BEHAVIORAL;