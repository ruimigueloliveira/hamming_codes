LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PARITY_BITS_CALCULATOR IS
  PORT( CODED_MESSAGE : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
		  PARITY_BIT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END PARITY_BITS_CALCULATOR;

ARCHITECTURE STRUCTURAL OF PARITY_BITS_CALCULATOR IS
BEGIN

	PARITY_BIT(0) <= CODED_MESSAGE(1-1) XOR CODED_MESSAGE(2-1)  XOR CODED_MESSAGE(3-1)  XOR CODED_MESSAGE(7-1)  XOR
						  CODED_MESSAGE(8-1) XOR CODED_MESSAGE(9-1)  XOR CODED_MESSAGE(11-1) XOR CODED_MESSAGE(12-1);
						  
	PARITY_BIT(1) <= CODED_MESSAGE(1-1) XOR CODED_MESSAGE(4-1)  XOR CODED_MESSAGE(5-1)  XOR CODED_MESSAGE(7-1)  XOR
						  CODED_MESSAGE(8-1) XOR CODED_MESSAGE(10-1) XOR CODED_MESSAGE(11-1) XOR CODED_MESSAGE(13-1);
						  
	PARITY_BIT(2) <= CODED_MESSAGE(2-1) XOR CODED_MESSAGE(4-1)  XOR CODED_MESSAGE(6-1)  XOR CODED_MESSAGE(7-1)  XOR
						  CODED_MESSAGE(9-1) XOR CODED_MESSAGE(10-1) XOR CODED_MESSAGE(11-1) XOR CODED_MESSAGE(14-1);
						  
	PARITY_BIT(3) <= CODED_MESSAGE(3-1) XOR CODED_MESSAGE(5-1)  XOR CODED_MESSAGE(6-1)  XOR CODED_MESSAGE(8-1)  XOR
						  CODED_MESSAGE(9-1) XOR CODED_MESSAGE(10-1) XOR CODED_MESSAGE(11-1) XOR CODED_MESSAGE(15-1);
						  
END STRUCTURAL;
