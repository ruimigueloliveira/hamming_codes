LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PARITY_BITS_CALCULATOR IS
  PORT( Y : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
		  PARITY_BIT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END PARITY_BITS_CALCULATOR;

ARCHITECTURE STRUCTURAL OF PARITY_BITS_CALCULATOR IS

-- LEVEL ONE
SIGNAL XOR_Y01_Y07, XOR_Y08_Y11, XOR_Y02_Y03, XOR_Y09_Y12, XOR_Y04_Y05, XOR_Y10_Y13, XOR_Y06_Y09, XOR_Y10_Y11, XOR_Y02_Y04, XOR_Y07_Y14, XOR_Y03_Y05, XOR_Y08_Y15: STD_LOGIC;

-- LEVEL TWO
SIGNAL XOR_Y01_Y07_Y08_Y11, XOR_Y02_Y03_Y09_Y12, XOR_Y04_Y05_Y10_Y13, XOR_Y06_Y09_Y10_Y11, XOR_Y02_Y04_Y07_Y14, XOR_Y03_Y05_Y08_Y15: STD_LOGIC;

BEGIN
	
	-- LEVEL ONE
	XOR_Y01_Y07 <= Y(0) XOR Y(6) ;
	XOR_Y08_Y11 <= Y(7) XOR Y(10);
	XOR_Y02_Y03 <= Y(1) XOR Y(2);
	XOR_Y09_Y12 <= Y(8) XOR Y(11);
	XOR_Y04_Y05 <= Y(3) XOR Y(4);
	XOR_Y10_Y13 <= Y(9) XOR Y(12);
	XOR_Y06_Y09 <= Y(5) XOR Y(8);
	XOR_Y10_Y11 <= Y(9) XOR Y(10);
	XOR_Y02_Y04 <= Y(1) XOR Y(3);
	XOR_Y07_Y14 <= Y(6) XOR Y(13);
	XOR_Y03_Y05 <= Y(2) XOR Y(4);
	XOR_Y08_Y15 <= Y(7) XOR Y(14);
	
	-- LEVEL TWO
	XOR_Y01_Y07_Y08_Y11 <= XOR_Y01_Y07 XOR XOR_Y08_Y11;
	XOR_Y02_Y03_Y09_Y12 <= XOR_Y02_Y03 XOR XOR_Y09_Y12;
	XOR_Y04_Y05_Y10_Y13 <= XOR_Y04_Y05 XOR XOR_Y10_Y13;
	XOR_Y06_Y09_Y10_Y11 <= XOR_Y06_Y09 XOR XOR_Y10_Y11;
	XOR_Y02_Y04_Y07_Y14 <= XOR_Y02_Y04 XOR XOR_Y07_Y14;
	XOR_Y03_Y05_Y08_Y15 <= XOR_Y03_Y05 XOR XOR_Y08_Y15;
	
	-- LEVEL THREE
	PARITY_BIT(0) <= XOR_Y01_Y07_Y08_Y11 XOR XOR_Y02_Y03_Y09_Y12; 
	PARITY_BIT(1) <= XOR_Y01_Y07_Y08_Y11 XOR XOR_Y04_Y05_Y10_Y13; 
	PARITY_BIT(2) <= XOR_Y06_Y09_Y10_Y11 XOR XOR_Y02_Y04_Y07_Y14; 
	PARITY_BIT(3) <= XOR_Y06_Y09_Y10_Y11 XOR XOR_Y03_Y05_Y08_Y15; 
						  
END STRUCTURAL;
