LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MULT4TO1 IS
	PORT (X00,X01,X10,X11: IN STD_LOGIC;
        S: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
        Y: OUT STD_LOGIC);
END MULT4TO1;

ARCHITECTURE BEHAVIORAL OF MULT4TO1 IS

SIGNAL M0OUT : STD_LOGIC;
SIGNAL M1OUT : STD_LOGIC;

BEGIN
	MULT0: WORK.MULT2TO1 PORT MAP (X00, X01, S(0), M0OUT);
	MULT1: WORK.MULT2TO1 PORT MAP (X10, X11, S(0), M1OUT);
	MULT2: WORK.MULT2TO1 PORT MAP (M0OUT, M1OUT, S(1), Y);
END BEHAVIORAL;