LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY AXORB IS
  PORT (A,B: IN STD_LOGIC;
        AXB: OUT STD_LOGIC);
END AXORB;

ARCHITECTURE STRUCTURAL OF AXORB IS
BEGIN
	AXB<=A XOR B;
END STRUCTURAL;

-----------------------------------------------

--LIBRARY IEEE;
--USE IEEE.STD_LOGIC_1164.ALL;
--
--ENTITY AORB IS
--  PORT (A,B: IN STD_LOGIC;
--        AAB: OUT STD_LOGIC);
--END AORB;
--
--ARCHITECTURE STRUCTURAL OF AORB IS
--BEGIN
--	AAB<=A OR B;
--END STRUCTURAL;

-----------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY NOTA IS
  PORT (A: IN STD_LOGIC;
        NA: OUT STD_LOGIC);
END NOTA;

ARCHITECTURE STRUCTURAL OF NOTA IS
BEGIN
	NA<=NOT A;
END STRUCTURAL;

-----------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY AANDB IS
  PORT (A,B: IN STD_LOGIC;
        AAB: OUT STD_LOGIC);
END AANDB;

ARCHITECTURE STRUCTURAL OF AANDB IS
BEGIN
	AAB<=A AND B;
END STRUCTURAL;

-----------------------------------------------

--FORNECIDO PELO PROFESSOR NO LROT_8BIT.VHD 
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MULT2TO1 IS
  PORT (X0, X1: IN STD_LOGIC;
        S: IN STD_LOGIC;
        Y: OUT STD_LOGIC);
END MULT2TO1;

ARCHITECTURE LOGICFUNCTION OF MULT2TO1 IS
BEGIN
  Y <= (X0 AND NOT S) OR (X1 AND S);
END LOGICFUNCTION;

-----------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MULT4TO1 IS
  PORT (X00,X01,X10,X11: IN STD_LOGIC;
        S: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
        Y: OUT STD_LOGIC);
END MULT4TO1;

ARCHITECTURE LOGICFUNCTION OF MULT4TO1 IS
SIGNAL M0OUT : STD_LOGIC;
SIGNAL M1OUT : STD_LOGIC;
BEGIN
	MULT0: WORK.MULT2TO1 PORT MAP (X00, X01, S(0), M0OUT);
	MULT1: WORK.MULT2TO1 PORT MAP (X10, X11, S(0), M1OUT);
	MULT2: WORK.MULT2TO1 PORT MAP (M0OUT, M1OUT, S(1), Y);
END LOGICFUNCTION;

-----------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY HALFADDER1BIT IS
  PORT (A,B : IN STD_LOGIC;
        S,COUT: OUT STD_LOGIC);
END HALFADDER1BIT;

ARCHITECTURE LOGICFUNCTION OF HALFADDER1BIT IS
SIGNAL S_XORAB : STD_LOGIC;
BEGIN
	XOR0: WORK.AXORB PORT MAP (A,B,S);
	AND0: WORK.AANDB PORT MAP (A,B,COUT);	
END LOGICFUNCTION;

-----------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY INC4BIT IS
  PORT (A : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        S : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		  OVERFLOW : OUT STD_LOGIC);
END INC4BIT;

ARCHITECTURE LOGICFUNCTION OF INC4BIT IS
SIGNAL S_COUT0 : STD_LOGIC;
SIGNAL S_COUT1 : STD_LOGIC;
SIGNAL S_COUT2 : STD_LOGIC;
BEGIN
	HA0: WORK.HALFADDER1BIT PORT MAP (A(0),'1',S(0),S_COUT0);
	HA1: WORK.HALFADDER1BIT PORT MAP (A(1),S_COUT0,S(1),S_COUT1);
	HA2: WORK.HALFADDER1BIT PORT MAP (A(2),S_COUT1,S(2),S_COUT2);
	HA3: WORK.HALFADDER1BIT PORT MAP (A(3),S_COUT2,S(3),OVERFLOW);
END LOGICFUNCTION;


-----------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY COUNTER4BIT IS
  PORT( CLK : IN STD_LOGIC;
		  NRST : IN STD_LOGIC;
		  CNT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		  OVERFLOW : OUT STD_LOGIC);
END COUNTER4BIT;

ARCHITECTURE STRUCTURAL OF COUNTER4BIT IS
SIGNAL S_REG : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL S_CNT : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN

	REG0 : WORK.FLIPFLOPDSIMUL PORT MAP (CLK,S_CNT(0),'1',NRST,S_REG(0),OPEN);
	REG1 : WORK.FLIPFLOPDSIMUL PORT MAP (CLK,S_CNT(1),'1',NRST,S_REG(1),OPEN);
	REG2 : WORK.FLIPFLOPDSIMUL PORT MAP (CLK,S_CNT(2),'1',NRST,S_REG(2),OPEN);
	REG3 : WORK.FLIPFLOPDSIMUL PORT MAP (CLK,S_CNT(3),'1',NRST,S_REG(3),OPEN);

	INC : WORK.INC4BIT PORT MAP (S_REG,S_CNT,OVERFLOW);
	CNT<=S_REG;
	
END STRUCTURAL;
