LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY CONTROL_UNIT IS
	PORT(ADDR: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		  CTRLBITS: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END CONTROL_UNIT;

ARCHITECTURE BEHAVIORAL OF CONTROL_UNIT IS

	TYPE TROM IS ARRAY (0 TO 14) OF STD_LOGIC_VECTOR(6 DOWNTO 0); 
	CONSTANT ROM_TABLE : TROM := (
		"1100000",
		"1010000",
		"1001000",
		"0110000",
		"0101000",
		"0011000",
		"1110000",
		"1101000",
		"1011000",
		"0111000",
		"1111000",
		"0000100",
		"0000101",
		"0000110",
		"0000111"
		);
		
BEGIN
		CTRLBITS <= ROM_TABLE(TO_INTEGER(UNSIGNED(ADDR)));
		
END BEHAVIORAL;